//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: LKB
// Engineer: Leonhard Neuhaus
// 
// Create Date: 27.11.2014 14:15:43
// Design Name: 
// Module Name: red_pitaya_iq_fgen_block
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//  
// This module outputs 4 signed signals: 
// sin(f*t), cos(f*t),sin(f*t+phi), cos(f*t+phi)
// The maximally positive signal is 2**(LUTBITS-1)-1
// The maximally negative signal is -(2**(LUTBITS-1)-1)
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
/*
###############################################################################
#    pyrpl - DSP servo controller for quantum optics with the RedPitaya
#    Copyright (C) 2014-2016  Leonhard Neuhaus  (neuhaus@spectro.jussieu.fr)
#
#    This program is free software: you can redistribute it and/or modify
#    it under the terms of the GNU General Public License as published by
#    the Free Software Foundation, either version 3 of the License, or
#    (at your option) any later version.
#
#    This program is distributed in the hope that it will be useful,
#    but WITHOUT ANY WARRANTY; without even the implied warranty of
#    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
#    GNU General Public License for more details.
#
#    You should have received a copy of the GNU General Public License
#    along with this program.  If not, see <http://www.gnu.org/licenses/>.
############################################################################### 
*/


module red_pitaya_iq_fgen_block #(
    parameter     LUTSZ     = 11,  
    parameter     LUTBITS   = 17,  
    parameter     PHASEBITS = 32 
)
(
    input clk_i,
    input rstn_i,
    input on,
    input sin_at_2f,
    input cos_at_2f,
    input sin_shifted_at_2f,
    input cos_shifted_at_2f,

    input  [PHASEBITS-1:0] start_phase,
    input  [PHASEBITS-1:0] shift_phase,
    output [LUTBITS-1:0] sin_o      ,
    output [LUTBITS-1:0] cos_o      ,
    output [LUTBITS-1:0] sin_shifted_o      ,
    output [LUTBITS-1:0] cos_shifted_o      ,
    output [PHASEBITS-1:0] phase_o // Output current phase - either of sin or sin_shifted
);

reg [LUTBITS-1:0] sin;
reg [LUTBITS-1:0] cos;
reg [LUTBITS-1:0] sin_shifted;
reg [LUTBITS-1:0] cos_shifted;
reg [PHASEBITS-1:0] phase_o_reg;

assign sin_o = sin;
assign sin_shifted_o = sin_shifted;
assign cos_o = cos;
assign cos_shifted_o = cos_shifted;

localparam QSHIFT = {{PHASEBITS-1{1'b0}},1'b1}  << (PHASEBITS-2);

//lut data block
reg [LUTBITS-1-1:0] lutrom [0:(1<<LUTSZ)-1];
reg [PHASEBITS-1:0] phase;

wire [PHASEBITS-1:0] wwphase1;
wire [PHASEBITS-1:0] wwphase2;
wire [PHASEBITS-1:0] wwphase3;
wire [PHASEBITS-1:0] wwphase4;
wire [LUTBITS-1:0] wphase1;
wire [LUTBITS-1:0] wphase2;
wire [LUTBITS-1:0] wphase3;
wire [LUTBITS-1:0] wphase4;
wire invertphase1;
wire invertphase2;
wire invertphase3;
wire invertphase4;
wire invertsignal1;
wire invertsignal2;
wire invertsignal3;
wire invertsignal4;
reg invertsignal1_reg;
reg invertsignal2_reg;
reg invertsignal3_reg;
reg invertsignal4_reg;
reg invertsignal1_reg_reg;
reg invertsignal2_reg_reg;
reg invertsignal3_reg_reg;
reg invertsignal4_reg_reg;
reg [LUTBITS-1:0] sin_reg;
reg [LUTBITS-1:0] cos_reg;
reg [LUTBITS-1:0] sin_shifted_reg;
reg [LUTBITS-1:0] cos_shifted_reg;

reg [LUTBITS-1:0] phase1;
reg [LUTBITS-1:0] phase2;
reg [LUTBITS-1:0] phase3;
reg [LUTBITS-1:0] phase4;

// in clock cycle n-1, phase is incremented (see far below in the else-block
// in clock cycle n,
//     - we assign wwphase1-4, the phase of the 4 subgenerators (possibly doubled phase counter for generation at 2f)
//     - we assign wphase1-4,
//     - we assign invertphase1-4, the flag telling if we are in the rising or falling quadrant of the sine
//     - we assign invertsignal1-4, the flag telling if we in the positive or negative sign of the sine

assign wwphase1 = sin_at_2f ? {phase[PHASEBITS-1:0],1'b0} : phase; // wwphase1 ready in cycle n
assign wwphase2 = cos_at_2f ? {phase[PHASEBITS-1:0],1'b0} + QSHIFT : phase + QSHIFT;
assign wwphase3 = sin_shifted_at_2f ? {phase[PHASEBITS-1:0],1'b0} + start_phase : phase + start_phase;
assign wwphase4 = cos_shifted_at_2f ? {phase[PHASEBITS-1:0],1'b0} + start_phase + QSHIFT : phase + start_phase + QSHIFT;
assign wphase1 = wwphase1[PHASEBITS-2-1:PHASEBITS-2-LUTSZ]; //wwphase1 ready in cycle n
assign wphase2 = wwphase2[PHASEBITS-2-1:PHASEBITS-2-LUTSZ];
assign wphase3 = wwphase3[PHASEBITS-2-1:PHASEBITS-2-LUTSZ];
assign wphase4 = wwphase4[PHASEBITS-2-1:PHASEBITS-2-LUTSZ];
assign invertphase1  = wwphase1[PHASEBITS-1-1];  //invertphase1 ready in cycle n
assign invertphase2  = wwphase2[PHASEBITS-1-1]; 
assign invertphase3  = wwphase3[PHASEBITS-1-1]; 
assign invertphase4  = wwphase4[PHASEBITS-1-1]; 
assign invertsignal1 = wwphase1[PHASEBITS-1]; //invertsignal1 ready in cycle n
assign invertsignal2 = wwphase2[PHASEBITS-1];
assign invertsignal3 = wwphase3[PHASEBITS-1];
assign invertsignal4 = wwphase4[PHASEBITS-1];

assign phase_o = phase_o_reg;

//main loop
always @(posedge clk_i) begin
    // 1) Next-phase computations:
    phase1 <= invertphase1 ? (~wphase1) : wphase1;  //phase1 ready in cycle n+1
    phase2 <= invertphase2 ? (~wphase2) : wphase2;
    phase3 <= invertphase3 ? (~wphase3) : wphase3;
    phase4 <= invertphase4 ? (~wphase4) : wphase4;

    // 2) Register the sign bits
    invertsignal1_reg <= invertsignal1; //invertsignal1_reg ready in cycle n+1
    invertsignal2_reg <= invertsignal2;
    invertsignal3_reg <= invertsignal3;
    invertsignal4_reg <= invertsignal4;
    invertsignal1_reg_reg <= invertsignal1_reg; //invertsignal1_reg_reg ready in cycle n+2
    invertsignal2_reg_reg <= invertsignal2_reg;
    invertsignal3_reg_reg <= invertsignal3_reg;
    invertsignal4_reg_reg <= invertsignal4_reg;

    // 3) Read LUT outputs for the next cycle
    sin_reg <= lutrom[phase1];    //sin_reg ready in cycle n+2
    cos_reg <= lutrom[phase2];
    sin_shifted_reg <= lutrom[phase3];
    cos_shifted_reg <= lutrom[phase4];

    // 4) Reset vs. Running State
    if (on==1'b0) begin // TODO: additional reset condition for syncing with ASG period possibly
        phase <= {PHASEBITS{1'b0}};
        phase_o_reg <= {PHASEBITS{1'b0}};
        sin <= {LUTBITS{1'b0}};
        cos <= {LUTBITS{1'b0}};
        sin_shifted <= {LUTBITS{1'b0}};
        cos_shifted <= {LUTBITS{1'b0}};
    end 
    else begin
        // 5) Advance the phase accumulator 
        phase <= phase + shift_phase; // new phase is ready in (arbitrary) cycle n

        // 6) Invert sign if needed
        sin <= invertsignal1_reg_reg ? ((~sin_reg)+'b1) : sin_reg;    //sin ready in cycle n+3  - based purely on signals that are ready in cycle n+2 -> timing correct, latency 3 cycles
        cos <= invertsignal2_reg_reg ? ((~cos_reg)+'b1) : cos_reg; 
        sin_shifted <= invertsignal3_reg_reg ? ((~sin_shifted_reg)+'b1) : sin_shifted_reg;  
        cos_shifted <= invertsignal4_reg_reg ? ((~cos_shifted_reg)+'b1) : cos_shifted_reg;
        phase_o_reg <= phase + shift_phase;  // TODO: maybe instead phase_o <= phase, schauen, wann welcher Wert ausgegeben sollte
    end
end

//LUT ROM
//created by this (unpolished) python code:
/*
LUTSZ = 11     #number of LUT entries
LUTBITS = 17   #LUT word size
def from_pyint(v,bitlength=14):
    v = int(v)
    if v < 0:
        v = v + 2**bitlength
    v= (v & (2**bitlength-1))
    return int(v)
data = np.zeros(2**LUTSZ,dtype=np.long)
for i in range(len(data)):
    data[i] = np.long(np.round((2**(LUTBITS-1)-1)*np.sin(((float(i)+0.5)/len(data))*0.5*np.pi)))
data = [from_pyint(v,bitlength=LUTBITS) for v in data]
plot(data)

print "reg [LUTBITS-1-1:0] lutrom [0:(1<<LUTSZ)-1];"
print ""
print "initial begin"
for i in range(len(data)):
    string = "   lutrom["+str(i)+"] = "+str(LUTBITS-1)+"'d"+str(data[i])+";"
    print string
print "end"
*/ 


initial begin
   lutrom[0] = 16'd25;
   lutrom[1] = 16'd75;
   lutrom[2] = 16'd126;
   lutrom[3] = 16'd176;
   lutrom[4] = 16'd226;
   lutrom[5] = 16'd276;
   lutrom[6] = 16'd327;
   lutrom[7] = 16'd377;
   lutrom[8] = 16'd427;
   lutrom[9] = 16'd478;
   lutrom[10] = 16'd528;
   lutrom[11] = 16'd578;
   lutrom[12] = 16'd628;
   lutrom[13] = 16'd679;
   lutrom[14] = 16'd729;
   lutrom[15] = 16'd779;
   lutrom[16] = 16'd829;
   lutrom[17] = 16'd880;
   lutrom[18] = 16'd930;
   lutrom[19] = 16'd980;
   lutrom[20] = 16'd1030;
   lutrom[21] = 16'd1081;
   lutrom[22] = 16'd1131;
   lutrom[23] = 16'd1181;
   lutrom[24] = 16'd1231;
   lutrom[25] = 16'd1282;
   lutrom[26] = 16'd1332;
   lutrom[27] = 16'd1382;
   lutrom[28] = 16'd1432;
   lutrom[29] = 16'd1483;
   lutrom[30] = 16'd1533;
   lutrom[31] = 16'd1583;
   lutrom[32] = 16'd1633;
   lutrom[33] = 16'd1684;
   lutrom[34] = 16'd1734;
   lutrom[35] = 16'd1784;
   lutrom[36] = 16'd1834;
   lutrom[37] = 16'd1885;
   lutrom[38] = 16'd1935;
   lutrom[39] = 16'd1985;
   lutrom[40] = 16'd2035;
   lutrom[41] = 16'd2086;
   lutrom[42] = 16'd2136;
   lutrom[43] = 16'd2186;
   lutrom[44] = 16'd2236;
   lutrom[45] = 16'd2287;
   lutrom[46] = 16'd2337;
   lutrom[47] = 16'd2387;
   lutrom[48] = 16'd2437;
   lutrom[49] = 16'd2488;
   lutrom[50] = 16'd2538;
   lutrom[51] = 16'd2588;
   lutrom[52] = 16'd2638;
   lutrom[53] = 16'd2688;
   lutrom[54] = 16'd2739;
   lutrom[55] = 16'd2789;
   lutrom[56] = 16'd2839;
   lutrom[57] = 16'd2889;
   lutrom[58] = 16'd2939;
   lutrom[59] = 16'd2990;
   lutrom[60] = 16'd3040;
   lutrom[61] = 16'd3090;
   lutrom[62] = 16'd3140;
   lutrom[63] = 16'd3191;
   lutrom[64] = 16'd3241;
   lutrom[65] = 16'd3291;
   lutrom[66] = 16'd3341;
   lutrom[67] = 16'd3391;
   lutrom[68] = 16'd3442;
   lutrom[69] = 16'd3492;
   lutrom[70] = 16'd3542;
   lutrom[71] = 16'd3592;
   lutrom[72] = 16'd3642;
   lutrom[73] = 16'd3693;
   lutrom[74] = 16'd3743;
   lutrom[75] = 16'd3793;
   lutrom[76] = 16'd3843;
   lutrom[77] = 16'd3893;
   lutrom[78] = 16'd3943;
   lutrom[79] = 16'd3994;
   lutrom[80] = 16'd4044;
   lutrom[81] = 16'd4094;
   lutrom[82] = 16'd4144;
   lutrom[83] = 16'd4194;
   lutrom[84] = 16'd4244;
   lutrom[85] = 16'd4295;
   lutrom[86] = 16'd4345;
   lutrom[87] = 16'd4395;
   lutrom[88] = 16'd4445;
   lutrom[89] = 16'd4495;
   lutrom[90] = 16'd4545;
   lutrom[91] = 16'd4595;
   lutrom[92] = 16'd4646;
   lutrom[93] = 16'd4696;
   lutrom[94] = 16'd4746;
   lutrom[95] = 16'd4796;
   lutrom[96] = 16'd4846;
   lutrom[97] = 16'd4896;
   lutrom[98] = 16'd4946;
   lutrom[99] = 16'd4996;
   lutrom[100] = 16'd5047;
   lutrom[101] = 16'd5097;
   lutrom[102] = 16'd5147;
   lutrom[103] = 16'd5197;
   lutrom[104] = 16'd5247;
   lutrom[105] = 16'd5297;
   lutrom[106] = 16'd5347;
   lutrom[107] = 16'd5397;
   lutrom[108] = 16'd5447;
   lutrom[109] = 16'd5498;
   lutrom[110] = 16'd5548;
   lutrom[111] = 16'd5598;
   lutrom[112] = 16'd5648;
   lutrom[113] = 16'd5698;
   lutrom[114] = 16'd5748;
   lutrom[115] = 16'd5798;
   lutrom[116] = 16'd5848;
   lutrom[117] = 16'd5898;
   lutrom[118] = 16'd5948;
   lutrom[119] = 16'd5998;
   lutrom[120] = 16'd6048;
   lutrom[121] = 16'd6098;
   lutrom[122] = 16'd6148;
   lutrom[123] = 16'd6198;
   lutrom[124] = 16'd6248;
   lutrom[125] = 16'd6298;
   lutrom[126] = 16'd6349;
   lutrom[127] = 16'd6399;
   lutrom[128] = 16'd6449;
   lutrom[129] = 16'd6499;
   lutrom[130] = 16'd6549;
   lutrom[131] = 16'd6599;
   lutrom[132] = 16'd6649;
   lutrom[133] = 16'd6699;
   lutrom[134] = 16'd6749;
   lutrom[135] = 16'd6799;
   lutrom[136] = 16'd6849;
   lutrom[137] = 16'd6899;
   lutrom[138] = 16'd6949;
   lutrom[139] = 16'd6999;
   lutrom[140] = 16'd7049;
   lutrom[141] = 16'd7099;
   lutrom[142] = 16'd7148;
   lutrom[143] = 16'd7198;
   lutrom[144] = 16'd7248;
   lutrom[145] = 16'd7298;
   lutrom[146] = 16'd7348;
   lutrom[147] = 16'd7398;
   lutrom[148] = 16'd7448;
   lutrom[149] = 16'd7498;
   lutrom[150] = 16'd7548;
   lutrom[151] = 16'd7598;
   lutrom[152] = 16'd7648;
   lutrom[153] = 16'd7698;
   lutrom[154] = 16'd7748;
   lutrom[155] = 16'd7798;
   lutrom[156] = 16'd7848;
   lutrom[157] = 16'd7897;
   lutrom[158] = 16'd7947;
   lutrom[159] = 16'd7997;
   lutrom[160] = 16'd8047;
   lutrom[161] = 16'd8097;
   lutrom[162] = 16'd8147;
   lutrom[163] = 16'd8197;
   lutrom[164] = 16'd8247;
   lutrom[165] = 16'd8296;
   lutrom[166] = 16'd8346;
   lutrom[167] = 16'd8396;
   lutrom[168] = 16'd8446;
   lutrom[169] = 16'd8496;
   lutrom[170] = 16'd8546;
   lutrom[171] = 16'd8596;
   lutrom[172] = 16'd8645;
   lutrom[173] = 16'd8695;
   lutrom[174] = 16'd8745;
   lutrom[175] = 16'd8795;
   lutrom[176] = 16'd8845;
   lutrom[177] = 16'd8894;
   lutrom[178] = 16'd8944;
   lutrom[179] = 16'd8994;
   lutrom[180] = 16'd9044;
   lutrom[181] = 16'd9094;
   lutrom[182] = 16'd9143;
   lutrom[183] = 16'd9193;
   lutrom[184] = 16'd9243;
   lutrom[185] = 16'd9293;
   lutrom[186] = 16'd9342;
   lutrom[187] = 16'd9392;
   lutrom[188] = 16'd9442;
   lutrom[189] = 16'd9492;
   lutrom[190] = 16'd9541;
   lutrom[191] = 16'd9591;
   lutrom[192] = 16'd9641;
   lutrom[193] = 16'd9691;
   lutrom[194] = 16'd9740;
   lutrom[195] = 16'd9790;
   lutrom[196] = 16'd9840;
   lutrom[197] = 16'd9889;
   lutrom[198] = 16'd9939;
   lutrom[199] = 16'd9989;
   lutrom[200] = 16'd10038;
   lutrom[201] = 16'd10088;
   lutrom[202] = 16'd10138;
   lutrom[203] = 16'd10187;
   lutrom[204] = 16'd10237;
   lutrom[205] = 16'd10287;
   lutrom[206] = 16'd10336;
   lutrom[207] = 16'd10386;
   lutrom[208] = 16'd10436;
   lutrom[209] = 16'd10485;
   lutrom[210] = 16'd10535;
   lutrom[211] = 16'd10584;
   lutrom[212] = 16'd10634;
   lutrom[213] = 16'd10684;
   lutrom[214] = 16'd10733;
   lutrom[215] = 16'd10783;
   lutrom[216] = 16'd10832;
   lutrom[217] = 16'd10882;
   lutrom[218] = 16'd10932;
   lutrom[219] = 16'd10981;
   lutrom[220] = 16'd11031;
   lutrom[221] = 16'd11080;
   lutrom[222] = 16'd11130;
   lutrom[223] = 16'd11179;
   lutrom[224] = 16'd11229;
   lutrom[225] = 16'd11278;
   lutrom[226] = 16'd11328;
   lutrom[227] = 16'd11377;
   lutrom[228] = 16'd11427;
   lutrom[229] = 16'd11476;
   lutrom[230] = 16'd11526;
   lutrom[231] = 16'd11575;
   lutrom[232] = 16'd11625;
   lutrom[233] = 16'd11674;
   lutrom[234] = 16'd11724;
   lutrom[235] = 16'd11773;
   lutrom[236] = 16'd11823;
   lutrom[237] = 16'd11872;
   lutrom[238] = 16'd11921;
   lutrom[239] = 16'd11971;
   lutrom[240] = 16'd12020;
   lutrom[241] = 16'd12070;
   lutrom[242] = 16'd12119;
   lutrom[243] = 16'd12168;
   lutrom[244] = 16'd12218;
   lutrom[245] = 16'd12267;
   lutrom[246] = 16'd12317;
   lutrom[247] = 16'd12366;
   lutrom[248] = 16'd12415;
   lutrom[249] = 16'd12465;
   lutrom[250] = 16'd12514;
   lutrom[251] = 16'd12563;
   lutrom[252] = 16'd12613;
   lutrom[253] = 16'd12662;
   lutrom[254] = 16'd12711;
   lutrom[255] = 16'd12761;
   lutrom[256] = 16'd12810;
   lutrom[257] = 16'd12859;
   lutrom[258] = 16'd12908;
   lutrom[259] = 16'd12958;
   lutrom[260] = 16'd13007;
   lutrom[261] = 16'd13056;
   lutrom[262] = 16'd13106;
   lutrom[263] = 16'd13155;
   lutrom[264] = 16'd13204;
   lutrom[265] = 16'd13253;
   lutrom[266] = 16'd13302;
   lutrom[267] = 16'd13352;
   lutrom[268] = 16'd13401;
   lutrom[269] = 16'd13450;
   lutrom[270] = 16'd13499;
   lutrom[271] = 16'd13548;
   lutrom[272] = 16'd13598;
   lutrom[273] = 16'd13647;
   lutrom[274] = 16'd13696;
   lutrom[275] = 16'd13745;
   lutrom[276] = 16'd13794;
   lutrom[277] = 16'd13843;
   lutrom[278] = 16'd13893;
   lutrom[279] = 16'd13942;
   lutrom[280] = 16'd13991;
   lutrom[281] = 16'd14040;
   lutrom[282] = 16'd14089;
   lutrom[283] = 16'd14138;
   lutrom[284] = 16'd14187;
   lutrom[285] = 16'd14236;
   lutrom[286] = 16'd14285;
   lutrom[287] = 16'd14334;
   lutrom[288] = 16'd14383;
   lutrom[289] = 16'd14432;
   lutrom[290] = 16'd14481;
   lutrom[291] = 16'd14530;
   lutrom[292] = 16'd14579;
   lutrom[293] = 16'd14628;
   lutrom[294] = 16'd14677;
   lutrom[295] = 16'd14726;
   lutrom[296] = 16'd14775;
   lutrom[297] = 16'd14824;
   lutrom[298] = 16'd14873;
   lutrom[299] = 16'd14922;
   lutrom[300] = 16'd14971;
   lutrom[301] = 16'd15020;
   lutrom[302] = 16'd15069;
   lutrom[303] = 16'd15118;
   lutrom[304] = 16'd15167;
   lutrom[305] = 16'd15216;
   lutrom[306] = 16'd15265;
   lutrom[307] = 16'd15314;
   lutrom[308] = 16'd15362;
   lutrom[309] = 16'd15411;
   lutrom[310] = 16'd15460;
   lutrom[311] = 16'd15509;
   lutrom[312] = 16'd15558;
   lutrom[313] = 16'd15607;
   lutrom[314] = 16'd15655;
   lutrom[315] = 16'd15704;
   lutrom[316] = 16'd15753;
   lutrom[317] = 16'd15802;
   lutrom[318] = 16'd15851;
   lutrom[319] = 16'd15899;
   lutrom[320] = 16'd15948;
   lutrom[321] = 16'd15997;
   lutrom[322] = 16'd16046;
   lutrom[323] = 16'd16094;
   lutrom[324] = 16'd16143;
   lutrom[325] = 16'd16192;
   lutrom[326] = 16'd16240;
   lutrom[327] = 16'd16289;
   lutrom[328] = 16'd16338;
   lutrom[329] = 16'd16386;
   lutrom[330] = 16'd16435;
   lutrom[331] = 16'd16484;
   lutrom[332] = 16'd16532;
   lutrom[333] = 16'd16581;
   lutrom[334] = 16'd16630;
   lutrom[335] = 16'd16678;
   lutrom[336] = 16'd16727;
   lutrom[337] = 16'd16776;
   lutrom[338] = 16'd16824;
   lutrom[339] = 16'd16873;
   lutrom[340] = 16'd16921;
   lutrom[341] = 16'd16970;
   lutrom[342] = 16'd17018;
   lutrom[343] = 16'd17067;
   lutrom[344] = 16'd17115;
   lutrom[345] = 16'd17164;
   lutrom[346] = 16'd17212;
   lutrom[347] = 16'd17261;
   lutrom[348] = 16'd17309;
   lutrom[349] = 16'd17358;
   lutrom[350] = 16'd17406;
   lutrom[351] = 16'd17455;
   lutrom[352] = 16'd17503;
   lutrom[353] = 16'd17552;
   lutrom[354] = 16'd17600;
   lutrom[355] = 16'd17649;
   lutrom[356] = 16'd17697;
   lutrom[357] = 16'd17745;
   lutrom[358] = 16'd17794;
   lutrom[359] = 16'd17842;
   lutrom[360] = 16'd17890;
   lutrom[361] = 16'd17939;
   lutrom[362] = 16'd17987;
   lutrom[363] = 16'd18035;
   lutrom[364] = 16'd18084;
   lutrom[365] = 16'd18132;
   lutrom[366] = 16'd18180;
   lutrom[367] = 16'd18229;
   lutrom[368] = 16'd18277;
   lutrom[369] = 16'd18325;
   lutrom[370] = 16'd18373;
   lutrom[371] = 16'd18422;
   lutrom[372] = 16'd18470;
   lutrom[373] = 16'd18518;
   lutrom[374] = 16'd18566;
   lutrom[375] = 16'd18615;
   lutrom[376] = 16'd18663;
   lutrom[377] = 16'd18711;
   lutrom[378] = 16'd18759;
   lutrom[379] = 16'd18807;
   lutrom[380] = 16'd18855;
   lutrom[381] = 16'd18904;
   lutrom[382] = 16'd18952;
   lutrom[383] = 16'd19000;
   lutrom[384] = 16'd19048;
   lutrom[385] = 16'd19096;
   lutrom[386] = 16'd19144;
   lutrom[387] = 16'd19192;
   lutrom[388] = 16'd19240;
   lutrom[389] = 16'd19288;
   lutrom[390] = 16'd19336;
   lutrom[391] = 16'd19384;
   lutrom[392] = 16'd19432;
   lutrom[393] = 16'd19480;
   lutrom[394] = 16'd19528;
   lutrom[395] = 16'd19576;
   lutrom[396] = 16'd19624;
   lutrom[397] = 16'd19672;
   lutrom[398] = 16'd19720;
   lutrom[399] = 16'd19768;
   lutrom[400] = 16'd19816;
   lutrom[401] = 16'd19864;
   lutrom[402] = 16'd19912;
   lutrom[403] = 16'd19960;
   lutrom[404] = 16'd20007;
   lutrom[405] = 16'd20055;
   lutrom[406] = 16'd20103;
   lutrom[407] = 16'd20151;
   lutrom[408] = 16'd20199;
   lutrom[409] = 16'd20247;
   lutrom[410] = 16'd20294;
   lutrom[411] = 16'd20342;
   lutrom[412] = 16'd20390;
   lutrom[413] = 16'd20438;
   lutrom[414] = 16'd20486;
   lutrom[415] = 16'd20533;
   lutrom[416] = 16'd20581;
   lutrom[417] = 16'd20629;
   lutrom[418] = 16'd20676;
   lutrom[419] = 16'd20724;
   lutrom[420] = 16'd20772;
   lutrom[421] = 16'd20819;
   lutrom[422] = 16'd20867;
   lutrom[423] = 16'd20915;
   lutrom[424] = 16'd20962;
   lutrom[425] = 16'd21010;
   lutrom[426] = 16'd21058;
   lutrom[427] = 16'd21105;
   lutrom[428] = 16'd21153;
   lutrom[429] = 16'd21200;
   lutrom[430] = 16'd21248;
   lutrom[431] = 16'd21295;
   lutrom[432] = 16'd21343;
   lutrom[433] = 16'd21390;
   lutrom[434] = 16'd21438;
   lutrom[435] = 16'd21485;
   lutrom[436] = 16'd21533;
   lutrom[437] = 16'd21580;
   lutrom[438] = 16'd21628;
   lutrom[439] = 16'd21675;
   lutrom[440] = 16'd21723;
   lutrom[441] = 16'd21770;
   lutrom[442] = 16'd21818;
   lutrom[443] = 16'd21865;
   lutrom[444] = 16'd21912;
   lutrom[445] = 16'd21960;
   lutrom[446] = 16'd22007;
   lutrom[447] = 16'd22054;
   lutrom[448] = 16'd22102;
   lutrom[449] = 16'd22149;
   lutrom[450] = 16'd22196;
   lutrom[451] = 16'd22244;
   lutrom[452] = 16'd22291;
   lutrom[453] = 16'd22338;
   lutrom[454] = 16'd22385;
   lutrom[455] = 16'd22433;
   lutrom[456] = 16'd22480;
   lutrom[457] = 16'd22527;
   lutrom[458] = 16'd22574;
   lutrom[459] = 16'd22621;
   lutrom[460] = 16'd22669;
   lutrom[461] = 16'd22716;
   lutrom[462] = 16'd22763;
   lutrom[463] = 16'd22810;
   lutrom[464] = 16'd22857;
   lutrom[465] = 16'd22904;
   lutrom[466] = 16'd22951;
   lutrom[467] = 16'd22998;
   lutrom[468] = 16'd23045;
   lutrom[469] = 16'd23093;
   lutrom[470] = 16'd23140;
   lutrom[471] = 16'd23187;
   lutrom[472] = 16'd23234;
   lutrom[473] = 16'd23281;
   lutrom[474] = 16'd23328;
   lutrom[475] = 16'd23375;
   lutrom[476] = 16'd23421;
   lutrom[477] = 16'd23468;
   lutrom[478] = 16'd23515;
   lutrom[479] = 16'd23562;
   lutrom[480] = 16'd23609;
   lutrom[481] = 16'd23656;
   lutrom[482] = 16'd23703;
   lutrom[483] = 16'd23750;
   lutrom[484] = 16'd23797;
   lutrom[485] = 16'd23843;
   lutrom[486] = 16'd23890;
   lutrom[487] = 16'd23937;
   lutrom[488] = 16'd23984;
   lutrom[489] = 16'd24031;
   lutrom[490] = 16'd24077;
   lutrom[491] = 16'd24124;
   lutrom[492] = 16'd24171;
   lutrom[493] = 16'd24218;
   lutrom[494] = 16'd24264;
   lutrom[495] = 16'd24311;
   lutrom[496] = 16'd24358;
   lutrom[497] = 16'd24404;
   lutrom[498] = 16'd24451;
   lutrom[499] = 16'd24498;
   lutrom[500] = 16'd24544;
   lutrom[501] = 16'd24591;
   lutrom[502] = 16'd24637;
   lutrom[503] = 16'd24684;
   lutrom[504] = 16'd24730;
   lutrom[505] = 16'd24777;
   lutrom[506] = 16'd24824;
   lutrom[507] = 16'd24870;
   lutrom[508] = 16'd24917;
   lutrom[509] = 16'd24963;
   lutrom[510] = 16'd25009;
   lutrom[511] = 16'd25056;
   lutrom[512] = 16'd25102;
   lutrom[513] = 16'd25149;
   lutrom[514] = 16'd25195;
   lutrom[515] = 16'd25242;
   lutrom[516] = 16'd25288;
   lutrom[517] = 16'd25334;
   lutrom[518] = 16'd25381;
   lutrom[519] = 16'd25427;
   lutrom[520] = 16'd25473;
   lutrom[521] = 16'd25520;
   lutrom[522] = 16'd25566;
   lutrom[523] = 16'd25612;
   lutrom[524] = 16'd25658;
   lutrom[525] = 16'd25705;
   lutrom[526] = 16'd25751;
   lutrom[527] = 16'd25797;
   lutrom[528] = 16'd25843;
   lutrom[529] = 16'd25890;
   lutrom[530] = 16'd25936;
   lutrom[531] = 16'd25982;
   lutrom[532] = 16'd26028;
   lutrom[533] = 16'd26074;
   lutrom[534] = 16'd26120;
   lutrom[535] = 16'd26166;
   lutrom[536] = 16'd26212;
   lutrom[537] = 16'd26258;
   lutrom[538] = 16'd26305;
   lutrom[539] = 16'd26351;
   lutrom[540] = 16'd26397;
   lutrom[541] = 16'd26443;
   lutrom[542] = 16'd26489;
   lutrom[543] = 16'd26535;
   lutrom[544] = 16'd26580;
   lutrom[545] = 16'd26626;
   lutrom[546] = 16'd26672;
   lutrom[547] = 16'd26718;
   lutrom[548] = 16'd26764;
   lutrom[549] = 16'd26810;
   lutrom[550] = 16'd26856;
   lutrom[551] = 16'd26902;
   lutrom[552] = 16'd26948;
   lutrom[553] = 16'd26993;
   lutrom[554] = 16'd27039;
   lutrom[555] = 16'd27085;
   lutrom[556] = 16'd27131;
   lutrom[557] = 16'd27176;
   lutrom[558] = 16'd27222;
   lutrom[559] = 16'd27268;
   lutrom[560] = 16'd27314;
   lutrom[561] = 16'd27359;
   lutrom[562] = 16'd27405;
   lutrom[563] = 16'd27451;
   lutrom[564] = 16'd27496;
   lutrom[565] = 16'd27542;
   lutrom[566] = 16'd27587;
   lutrom[567] = 16'd27633;
   lutrom[568] = 16'd27679;
   lutrom[569] = 16'd27724;
   lutrom[570] = 16'd27770;
   lutrom[571] = 16'd27815;
   lutrom[572] = 16'd27861;
   lutrom[573] = 16'd27906;
   lutrom[574] = 16'd27952;
   lutrom[575] = 16'd27997;
   lutrom[576] = 16'd28043;
   lutrom[577] = 16'd28088;
   lutrom[578] = 16'd28133;
   lutrom[579] = 16'd28179;
   lutrom[580] = 16'd28224;
   lutrom[581] = 16'd28269;
   lutrom[582] = 16'd28315;
   lutrom[583] = 16'd28360;
   lutrom[584] = 16'd28405;
   lutrom[585] = 16'd28451;
   lutrom[586] = 16'd28496;
   lutrom[587] = 16'd28541;
   lutrom[588] = 16'd28587;
   lutrom[589] = 16'd28632;
   lutrom[590] = 16'd28677;
   lutrom[591] = 16'd28722;
   lutrom[592] = 16'd28767;
   lutrom[593] = 16'd28812;
   lutrom[594] = 16'd28858;
   lutrom[595] = 16'd28903;
   lutrom[596] = 16'd28948;
   lutrom[597] = 16'd28993;
   lutrom[598] = 16'd29038;
   lutrom[599] = 16'd29083;
   lutrom[600] = 16'd29128;
   lutrom[601] = 16'd29173;
   lutrom[602] = 16'd29218;
   lutrom[603] = 16'd29263;
   lutrom[604] = 16'd29308;
   lutrom[605] = 16'd29353;
   lutrom[606] = 16'd29398;
   lutrom[607] = 16'd29443;
   lutrom[608] = 16'd29488;
   lutrom[609] = 16'd29533;
   lutrom[610] = 16'd29577;
   lutrom[611] = 16'd29622;
   lutrom[612] = 16'd29667;
   lutrom[613] = 16'd29712;
   lutrom[614] = 16'd29757;
   lutrom[615] = 16'd29802;
   lutrom[616] = 16'd29846;
   lutrom[617] = 16'd29891;
   lutrom[618] = 16'd29936;
   lutrom[619] = 16'd29980;
   lutrom[620] = 16'd30025;
   lutrom[621] = 16'd30070;
   lutrom[622] = 16'd30114;
   lutrom[623] = 16'd30159;
   lutrom[624] = 16'd30204;
   lutrom[625] = 16'd30248;
   lutrom[626] = 16'd30293;
   lutrom[627] = 16'd30337;
   lutrom[628] = 16'd30382;
   lutrom[629] = 16'd30427;
   lutrom[630] = 16'd30471;
   lutrom[631] = 16'd30516;
   lutrom[632] = 16'd30560;
   lutrom[633] = 16'd30604;
   lutrom[634] = 16'd30649;
   lutrom[635] = 16'd30693;
   lutrom[636] = 16'd30738;
   lutrom[637] = 16'd30782;
   lutrom[638] = 16'd30826;
   lutrom[639] = 16'd30871;
   lutrom[640] = 16'd30915;
   lutrom[641] = 16'd30959;
   lutrom[642] = 16'd31004;
   lutrom[643] = 16'd31048;
   lutrom[644] = 16'd31092;
   lutrom[645] = 16'd31137;
   lutrom[646] = 16'd31181;
   lutrom[647] = 16'd31225;
   lutrom[648] = 16'd31269;
   lutrom[649] = 16'd31313;
   lutrom[650] = 16'd31357;
   lutrom[651] = 16'd31402;
   lutrom[652] = 16'd31446;
   lutrom[653] = 16'd31490;
   lutrom[654] = 16'd31534;
   lutrom[655] = 16'd31578;
   lutrom[656] = 16'd31622;
   lutrom[657] = 16'd31666;
   lutrom[658] = 16'd31710;
   lutrom[659] = 16'd31754;
   lutrom[660] = 16'd31798;
   lutrom[661] = 16'd31842;
   lutrom[662] = 16'd31886;
   lutrom[663] = 16'd31930;
   lutrom[664] = 16'd31974;
   lutrom[665] = 16'd32017;
   lutrom[666] = 16'd32061;
   lutrom[667] = 16'd32105;
   lutrom[668] = 16'd32149;
   lutrom[669] = 16'd32193;
   lutrom[670] = 16'd32236;
   lutrom[671] = 16'd32280;
   lutrom[672] = 16'd32324;
   lutrom[673] = 16'd32368;
   lutrom[674] = 16'd32411;
   lutrom[675] = 16'd32455;
   lutrom[676] = 16'd32499;
   lutrom[677] = 16'd32542;
   lutrom[678] = 16'd32586;
   lutrom[679] = 16'd32630;
   lutrom[680] = 16'd32673;
   lutrom[681] = 16'd32717;
   lutrom[682] = 16'd32760;
   lutrom[683] = 16'd32804;
   lutrom[684] = 16'd32847;
   lutrom[685] = 16'd32891;
   lutrom[686] = 16'd32934;
   lutrom[687] = 16'd32978;
   lutrom[688] = 16'd33021;
   lutrom[689] = 16'd33065;
   lutrom[690] = 16'd33108;
   lutrom[691] = 16'd33151;
   lutrom[692] = 16'd33195;
   lutrom[693] = 16'd33238;
   lutrom[694] = 16'd33281;
   lutrom[695] = 16'd33325;
   lutrom[696] = 16'd33368;
   lutrom[697] = 16'd33411;
   lutrom[698] = 16'd33454;
   lutrom[699] = 16'd33498;
   lutrom[700] = 16'd33541;
   lutrom[701] = 16'd33584;
   lutrom[702] = 16'd33627;
   lutrom[703] = 16'd33670;
   lutrom[704] = 16'd33713;
   lutrom[705] = 16'd33756;
   lutrom[706] = 16'd33799;
   lutrom[707] = 16'd33842;
   lutrom[708] = 16'd33886;
   lutrom[709] = 16'd33929;
   lutrom[710] = 16'd33972;
   lutrom[711] = 16'd34015;
   lutrom[712] = 16'd34057;
   lutrom[713] = 16'd34100;
   lutrom[714] = 16'd34143;
   lutrom[715] = 16'd34186;
   lutrom[716] = 16'd34229;
   lutrom[717] = 16'd34272;
   lutrom[718] = 16'd34315;
   lutrom[719] = 16'd34358;
   lutrom[720] = 16'd34400;
   lutrom[721] = 16'd34443;
   lutrom[722] = 16'd34486;
   lutrom[723] = 16'd34529;
   lutrom[724] = 16'd34571;
   lutrom[725] = 16'd34614;
   lutrom[726] = 16'd34657;
   lutrom[727] = 16'd34699;
   lutrom[728] = 16'd34742;
   lutrom[729] = 16'd34785;
   lutrom[730] = 16'd34827;
   lutrom[731] = 16'd34870;
   lutrom[732] = 16'd34912;
   lutrom[733] = 16'd34955;
   lutrom[734] = 16'd34997;
   lutrom[735] = 16'd35040;
   lutrom[736] = 16'd35082;
   lutrom[737] = 16'd35125;
   lutrom[738] = 16'd35167;
   lutrom[739] = 16'd35210;
   lutrom[740] = 16'd35252;
   lutrom[741] = 16'd35294;
   lutrom[742] = 16'd35337;
   lutrom[743] = 16'd35379;
   lutrom[744] = 16'd35421;
   lutrom[745] = 16'd35464;
   lutrom[746] = 16'd35506;
   lutrom[747] = 16'd35548;
   lutrom[748] = 16'd35590;
   lutrom[749] = 16'd35632;
   lutrom[750] = 16'd35675;
   lutrom[751] = 16'd35717;
   lutrom[752] = 16'd35759;
   lutrom[753] = 16'd35801;
   lutrom[754] = 16'd35843;
   lutrom[755] = 16'd35885;
   lutrom[756] = 16'd35927;
   lutrom[757] = 16'd35969;
   lutrom[758] = 16'd36011;
   lutrom[759] = 16'd36053;
   lutrom[760] = 16'd36095;
   lutrom[761] = 16'd36137;
   lutrom[762] = 16'd36179;
   lutrom[763] = 16'd36221;
   lutrom[764] = 16'd36263;
   lutrom[765] = 16'd36305;
   lutrom[766] = 16'd36347;
   lutrom[767] = 16'd36388;
   lutrom[768] = 16'd36430;
   lutrom[769] = 16'd36472;
   lutrom[770] = 16'd36514;
   lutrom[771] = 16'd36555;
   lutrom[772] = 16'd36597;
   lutrom[773] = 16'd36639;
   lutrom[774] = 16'd36680;
   lutrom[775] = 16'd36722;
   lutrom[776] = 16'd36764;
   lutrom[777] = 16'd36805;
   lutrom[778] = 16'd36847;
   lutrom[779] = 16'd36888;
   lutrom[780] = 16'd36930;
   lutrom[781] = 16'd36972;
   lutrom[782] = 16'd37013;
   lutrom[783] = 16'd37055;
   lutrom[784] = 16'd37096;
   lutrom[785] = 16'd37137;
   lutrom[786] = 16'd37179;
   lutrom[787] = 16'd37220;
   lutrom[788] = 16'd37262;
   lutrom[789] = 16'd37303;
   lutrom[790] = 16'd37344;
   lutrom[791] = 16'd37385;
   lutrom[792] = 16'd37427;
   lutrom[793] = 16'd37468;
   lutrom[794] = 16'd37509;
   lutrom[795] = 16'd37550;
   lutrom[796] = 16'd37592;
   lutrom[797] = 16'd37633;
   lutrom[798] = 16'd37674;
   lutrom[799] = 16'd37715;
   lutrom[800] = 16'd37756;
   lutrom[801] = 16'd37797;
   lutrom[802] = 16'd37838;
   lutrom[803] = 16'd37879;
   lutrom[804] = 16'd37920;
   lutrom[805] = 16'd37961;
   lutrom[806] = 16'd38002;
   lutrom[807] = 16'd38043;
   lutrom[808] = 16'd38084;
   lutrom[809] = 16'd38125;
   lutrom[810] = 16'd38166;
   lutrom[811] = 16'd38207;
   lutrom[812] = 16'd38248;
   lutrom[813] = 16'd38288;
   lutrom[814] = 16'd38329;
   lutrom[815] = 16'd38370;
   lutrom[816] = 16'd38411;
   lutrom[817] = 16'd38451;
   lutrom[818] = 16'd38492;
   lutrom[819] = 16'd38533;
   lutrom[820] = 16'd38573;
   lutrom[821] = 16'd38614;
   lutrom[822] = 16'd38655;
   lutrom[823] = 16'd38695;
   lutrom[824] = 16'd38736;
   lutrom[825] = 16'd38776;
   lutrom[826] = 16'd38817;
   lutrom[827] = 16'd38857;
   lutrom[828] = 16'd38898;
   lutrom[829] = 16'd38938;
   lutrom[830] = 16'd38979;
   lutrom[831] = 16'd39019;
   lutrom[832] = 16'd39059;
   lutrom[833] = 16'd39100;
   lutrom[834] = 16'd39140;
   lutrom[835] = 16'd39180;
   lutrom[836] = 16'd39221;
   lutrom[837] = 16'd39261;
   lutrom[838] = 16'd39301;
   lutrom[839] = 16'd39341;
   lutrom[840] = 16'd39381;
   lutrom[841] = 16'd39422;
   lutrom[842] = 16'd39462;
   lutrom[843] = 16'd39502;
   lutrom[844] = 16'd39542;
   lutrom[845] = 16'd39582;
   lutrom[846] = 16'd39622;
   lutrom[847] = 16'd39662;
   lutrom[848] = 16'd39702;
   lutrom[849] = 16'd39742;
   lutrom[850] = 16'd39782;
   lutrom[851] = 16'd39822;
   lutrom[852] = 16'd39862;
   lutrom[853] = 16'd39902;
   lutrom[854] = 16'd39942;
   lutrom[855] = 16'd39982;
   lutrom[856] = 16'd40021;
   lutrom[857] = 16'd40061;
   lutrom[858] = 16'd40101;
   lutrom[859] = 16'd40141;
   lutrom[860] = 16'd40180;
   lutrom[861] = 16'd40220;
   lutrom[862] = 16'd40260;
   lutrom[863] = 16'd40299;
   lutrom[864] = 16'd40339;
   lutrom[865] = 16'd40379;
   lutrom[866] = 16'd40418;
   lutrom[867] = 16'd40458;
   lutrom[868] = 16'd40497;
   lutrom[869] = 16'd40537;
   lutrom[870] = 16'd40576;
   lutrom[871] = 16'd40616;
   lutrom[872] = 16'd40655;
   lutrom[873] = 16'd40695;
   lutrom[874] = 16'd40734;
   lutrom[875] = 16'd40773;
   lutrom[876] = 16'd40813;
   lutrom[877] = 16'd40852;
   lutrom[878] = 16'd40891;
   lutrom[879] = 16'd40931;
   lutrom[880] = 16'd40970;
   lutrom[881] = 16'd41009;
   lutrom[882] = 16'd41048;
   lutrom[883] = 16'd41087;
   lutrom[884] = 16'd41127;
   lutrom[885] = 16'd41166;
   lutrom[886] = 16'd41205;
   lutrom[887] = 16'd41244;
   lutrom[888] = 16'd41283;
   lutrom[889] = 16'd41322;
   lutrom[890] = 16'd41361;
   lutrom[891] = 16'd41400;
   lutrom[892] = 16'd41439;
   lutrom[893] = 16'd41478;
   lutrom[894] = 16'd41517;
   lutrom[895] = 16'd41556;
   lutrom[896] = 16'd41594;
   lutrom[897] = 16'd41633;
   lutrom[898] = 16'd41672;
   lutrom[899] = 16'd41711;
   lutrom[900] = 16'd41750;
   lutrom[901] = 16'd41788;
   lutrom[902] = 16'd41827;
   lutrom[903] = 16'd41866;
   lutrom[904] = 16'd41904;
   lutrom[905] = 16'd41943;
   lutrom[906] = 16'd41982;
   lutrom[907] = 16'd42020;
   lutrom[908] = 16'd42059;
   lutrom[909] = 16'd42097;
   lutrom[910] = 16'd42136;
   lutrom[911] = 16'd42174;
   lutrom[912] = 16'd42213;
   lutrom[913] = 16'd42251;
   lutrom[914] = 16'd42290;
   lutrom[915] = 16'd42328;
   lutrom[916] = 16'd42366;
   lutrom[917] = 16'd42405;
   lutrom[918] = 16'd42443;
   lutrom[919] = 16'd42481;
   lutrom[920] = 16'd42520;
   lutrom[921] = 16'd42558;
   lutrom[922] = 16'd42596;
   lutrom[923] = 16'd42634;
   lutrom[924] = 16'd42672;
   lutrom[925] = 16'd42710;
   lutrom[926] = 16'd42749;
   lutrom[927] = 16'd42787;
   lutrom[928] = 16'd42825;
   lutrom[929] = 16'd42863;
   lutrom[930] = 16'd42901;
   lutrom[931] = 16'd42939;
   lutrom[932] = 16'd42977;
   lutrom[933] = 16'd43015;
   lutrom[934] = 16'd43053;
   lutrom[935] = 16'd43090;
   lutrom[936] = 16'd43128;
   lutrom[937] = 16'd43166;
   lutrom[938] = 16'd43204;
   lutrom[939] = 16'd43242;
   lutrom[940] = 16'd43279;
   lutrom[941] = 16'd43317;
   lutrom[942] = 16'd43355;
   lutrom[943] = 16'd43393;
   lutrom[944] = 16'd43430;
   lutrom[945] = 16'd43468;
   lutrom[946] = 16'd43505;
   lutrom[947] = 16'd43543;
   lutrom[948] = 16'd43581;
   lutrom[949] = 16'd43618;
   lutrom[950] = 16'd43656;
   lutrom[951] = 16'd43693;
   lutrom[952] = 16'd43731;
   lutrom[953] = 16'd43768;
   lutrom[954] = 16'd43805;
   lutrom[955] = 16'd43843;
   lutrom[956] = 16'd43880;
   lutrom[957] = 16'd43917;
   lutrom[958] = 16'd43955;
   lutrom[959] = 16'd43992;
   lutrom[960] = 16'd44029;
   lutrom[961] = 16'd44066;
   lutrom[962] = 16'd44104;
   lutrom[963] = 16'd44141;
   lutrom[964] = 16'd44178;
   lutrom[965] = 16'd44215;
   lutrom[966] = 16'd44252;
   lutrom[967] = 16'd44289;
   lutrom[968] = 16'd44326;
   lutrom[969] = 16'd44363;
   lutrom[970] = 16'd44400;
   lutrom[971] = 16'd44437;
   lutrom[972] = 16'd44474;
   lutrom[973] = 16'd44511;
   lutrom[974] = 16'd44548;
   lutrom[975] = 16'd44585;
   lutrom[976] = 16'd44622;
   lutrom[977] = 16'd44658;
   lutrom[978] = 16'd44695;
   lutrom[979] = 16'd44732;
   lutrom[980] = 16'd44769;
   lutrom[981] = 16'd44805;
   lutrom[982] = 16'd44842;
   lutrom[983] = 16'd44879;
   lutrom[984] = 16'd44915;
   lutrom[985] = 16'd44952;
   lutrom[986] = 16'd44988;
   lutrom[987] = 16'd45025;
   lutrom[988] = 16'd45061;
   lutrom[989] = 16'd45098;
   lutrom[990] = 16'd45134;
   lutrom[991] = 16'd45171;
   lutrom[992] = 16'd45207;
   lutrom[993] = 16'd45244;
   lutrom[994] = 16'd45280;
   lutrom[995] = 16'd45316;
   lutrom[996] = 16'd45353;
   lutrom[997] = 16'd45389;
   lutrom[998] = 16'd45425;
   lutrom[999] = 16'd45461;
   lutrom[1000] = 16'd45498;
   lutrom[1001] = 16'd45534;
   lutrom[1002] = 16'd45570;
   lutrom[1003] = 16'd45606;
   lutrom[1004] = 16'd45642;
   lutrom[1005] = 16'd45678;
   lutrom[1006] = 16'd45714;
   lutrom[1007] = 16'd45750;
   lutrom[1008] = 16'd45786;
   lutrom[1009] = 16'd45822;
   lutrom[1010] = 16'd45858;
   lutrom[1011] = 16'd45894;
   lutrom[1012] = 16'd45930;
   lutrom[1013] = 16'd45966;
   lutrom[1014] = 16'd46001;
   lutrom[1015] = 16'd46037;
   lutrom[1016] = 16'd46073;
   lutrom[1017] = 16'd46109;
   lutrom[1018] = 16'd46144;
   lutrom[1019] = 16'd46180;
   lutrom[1020] = 16'd46216;
   lutrom[1021] = 16'd46251;
   lutrom[1022] = 16'd46287;
   lutrom[1023] = 16'd46322;
   lutrom[1024] = 16'd46358;
   lutrom[1025] = 16'd46394;
   lutrom[1026] = 16'd46429;
   lutrom[1027] = 16'd46464;
   lutrom[1028] = 16'd46500;
   lutrom[1029] = 16'd46535;
   lutrom[1030] = 16'd46571;
   lutrom[1031] = 16'd46606;
   lutrom[1032] = 16'd46641;
   lutrom[1033] = 16'd46677;
   lutrom[1034] = 16'd46712;
   lutrom[1035] = 16'd46747;
   lutrom[1036] = 16'd46782;
   lutrom[1037] = 16'd46818;
   lutrom[1038] = 16'd46853;
   lutrom[1039] = 16'd46888;
   lutrom[1040] = 16'd46923;
   lutrom[1041] = 16'd46958;
   lutrom[1042] = 16'd46993;
   lutrom[1043] = 16'd47028;
   lutrom[1044] = 16'd47063;
   lutrom[1045] = 16'd47098;
   lutrom[1046] = 16'd47133;
   lutrom[1047] = 16'd47168;
   lutrom[1048] = 16'd47203;
   lutrom[1049] = 16'd47238;
   lutrom[1050] = 16'd47272;
   lutrom[1051] = 16'd47307;
   lutrom[1052] = 16'd47342;
   lutrom[1053] = 16'd47377;
   lutrom[1054] = 16'd47412;
   lutrom[1055] = 16'd47446;
   lutrom[1056] = 16'd47481;
   lutrom[1057] = 16'd47515;
   lutrom[1058] = 16'd47550;
   lutrom[1059] = 16'd47585;
   lutrom[1060] = 16'd47619;
   lutrom[1061] = 16'd47654;
   lutrom[1062] = 16'd47688;
   lutrom[1063] = 16'd47723;
   lutrom[1064] = 16'd47757;
   lutrom[1065] = 16'd47792;
   lutrom[1066] = 16'd47826;
   lutrom[1067] = 16'd47860;
   lutrom[1068] = 16'd47895;
   lutrom[1069] = 16'd47929;
   lutrom[1070] = 16'd47963;
   lutrom[1071] = 16'd47997;
   lutrom[1072] = 16'd48032;
   lutrom[1073] = 16'd48066;
   lutrom[1074] = 16'd48100;
   lutrom[1075] = 16'd48134;
   lutrom[1076] = 16'd48168;
   lutrom[1077] = 16'd48202;
   lutrom[1078] = 16'd48236;
   lutrom[1079] = 16'd48270;
   lutrom[1080] = 16'd48304;
   lutrom[1081] = 16'd48338;
   lutrom[1082] = 16'd48372;
   lutrom[1083] = 16'd48406;
   lutrom[1084] = 16'd48440;
   lutrom[1085] = 16'd48474;
   lutrom[1086] = 16'd48508;
   lutrom[1087] = 16'd48541;
   lutrom[1088] = 16'd48575;
   lutrom[1089] = 16'd48609;
   lutrom[1090] = 16'd48643;
   lutrom[1091] = 16'd48676;
   lutrom[1092] = 16'd48710;
   lutrom[1093] = 16'd48743;
   lutrom[1094] = 16'd48777;
   lutrom[1095] = 16'd48811;
   lutrom[1096] = 16'd48844;
   lutrom[1097] = 16'd48878;
   lutrom[1098] = 16'd48911;
   lutrom[1099] = 16'd48945;
   lutrom[1100] = 16'd48978;
   lutrom[1101] = 16'd49011;
   lutrom[1102] = 16'd49045;
   lutrom[1103] = 16'd49078;
   lutrom[1104] = 16'd49111;
   lutrom[1105] = 16'd49145;
   lutrom[1106] = 16'd49178;
   lutrom[1107] = 16'd49211;
   lutrom[1108] = 16'd49244;
   lutrom[1109] = 16'd49277;
   lutrom[1110] = 16'd49310;
   lutrom[1111] = 16'd49344;
   lutrom[1112] = 16'd49377;
   lutrom[1113] = 16'd49410;
   lutrom[1114] = 16'd49443;
   lutrom[1115] = 16'd49476;
   lutrom[1116] = 16'd49509;
   lutrom[1117] = 16'd49542;
   lutrom[1118] = 16'd49574;
   lutrom[1119] = 16'd49607;
   lutrom[1120] = 16'd49640;
   lutrom[1121] = 16'd49673;
   lutrom[1122] = 16'd49706;
   lutrom[1123] = 16'd49738;
   lutrom[1124] = 16'd49771;
   lutrom[1125] = 16'd49804;
   lutrom[1126] = 16'd49836;
   lutrom[1127] = 16'd49869;
   lutrom[1128] = 16'd49902;
   lutrom[1129] = 16'd49934;
   lutrom[1130] = 16'd49967;
   lutrom[1131] = 16'd49999;
   lutrom[1132] = 16'd50032;
   lutrom[1133] = 16'd50064;
   lutrom[1134] = 16'd50097;
   lutrom[1135] = 16'd50129;
   lutrom[1136] = 16'd50161;
   lutrom[1137] = 16'd50194;
   lutrom[1138] = 16'd50226;
   lutrom[1139] = 16'd50258;
   lutrom[1140] = 16'd50291;
   lutrom[1141] = 16'd50323;
   lutrom[1142] = 16'd50355;
   lutrom[1143] = 16'd50387;
   lutrom[1144] = 16'd50419;
   lutrom[1145] = 16'd50451;
   lutrom[1146] = 16'd50483;
   lutrom[1147] = 16'd50515;
   lutrom[1148] = 16'd50547;
   lutrom[1149] = 16'd50579;
   lutrom[1150] = 16'd50611;
   lutrom[1151] = 16'd50643;
   lutrom[1152] = 16'd50675;
   lutrom[1153] = 16'd50707;
   lutrom[1154] = 16'd50739;
   lutrom[1155] = 16'd50771;
   lutrom[1156] = 16'd50802;
   lutrom[1157] = 16'd50834;
   lutrom[1158] = 16'd50866;
   lutrom[1159] = 16'd50898;
   lutrom[1160] = 16'd50929;
   lutrom[1161] = 16'd50961;
   lutrom[1162] = 16'd50992;
   lutrom[1163] = 16'd51024;
   lutrom[1164] = 16'd51056;
   lutrom[1165] = 16'd51087;
   lutrom[1166] = 16'd51118;
   lutrom[1167] = 16'd51150;
   lutrom[1168] = 16'd51181;
   lutrom[1169] = 16'd51213;
   lutrom[1170] = 16'd51244;
   lutrom[1171] = 16'd51275;
   lutrom[1172] = 16'd51307;
   lutrom[1173] = 16'd51338;
   lutrom[1174] = 16'd51369;
   lutrom[1175] = 16'd51400;
   lutrom[1176] = 16'd51431;
   lutrom[1177] = 16'd51463;
   lutrom[1178] = 16'd51494;
   lutrom[1179] = 16'd51525;
   lutrom[1180] = 16'd51556;
   lutrom[1181] = 16'd51587;
   lutrom[1182] = 16'd51618;
   lutrom[1183] = 16'd51649;
   lutrom[1184] = 16'd51680;
   lutrom[1185] = 16'd51711;
   lutrom[1186] = 16'd51741;
   lutrom[1187] = 16'd51772;
   lutrom[1188] = 16'd51803;
   lutrom[1189] = 16'd51834;
   lutrom[1190] = 16'd51865;
   lutrom[1191] = 16'd51895;
   lutrom[1192] = 16'd51926;
   lutrom[1193] = 16'd51957;
   lutrom[1194] = 16'd51987;
   lutrom[1195] = 16'd52018;
   lutrom[1196] = 16'd52048;
   lutrom[1197] = 16'd52079;
   lutrom[1198] = 16'd52109;
   lutrom[1199] = 16'd52140;
   lutrom[1200] = 16'd52170;
   lutrom[1201] = 16'd52201;
   lutrom[1202] = 16'd52231;
   lutrom[1203] = 16'd52262;
   lutrom[1204] = 16'd52292;
   lutrom[1205] = 16'd52322;
   lutrom[1206] = 16'd52352;
   lutrom[1207] = 16'd52383;
   lutrom[1208] = 16'd52413;
   lutrom[1209] = 16'd52443;
   lutrom[1210] = 16'd52473;
   lutrom[1211] = 16'd52503;
   lutrom[1212] = 16'd52533;
   lutrom[1213] = 16'd52563;
   lutrom[1214] = 16'd52593;
   lutrom[1215] = 16'd52623;
   lutrom[1216] = 16'd52653;
   lutrom[1217] = 16'd52683;
   lutrom[1218] = 16'd52713;
   lutrom[1219] = 16'd52743;
   lutrom[1220] = 16'd52773;
   lutrom[1221] = 16'd52802;
   lutrom[1222] = 16'd52832;
   lutrom[1223] = 16'd52862;
   lutrom[1224] = 16'd52892;
   lutrom[1225] = 16'd52921;
   lutrom[1226] = 16'd52951;
   lutrom[1227] = 16'd52980;
   lutrom[1228] = 16'd53010;
   lutrom[1229] = 16'd53040;
   lutrom[1230] = 16'd53069;
   lutrom[1231] = 16'd53099;
   lutrom[1232] = 16'd53128;
   lutrom[1233] = 16'd53157;
   lutrom[1234] = 16'd53187;
   lutrom[1235] = 16'd53216;
   lutrom[1236] = 16'd53245;
   lutrom[1237] = 16'd53275;
   lutrom[1238] = 16'd53304;
   lutrom[1239] = 16'd53333;
   lutrom[1240] = 16'd53362;
   lutrom[1241] = 16'd53392;
   lutrom[1242] = 16'd53421;
   lutrom[1243] = 16'd53450;
   lutrom[1244] = 16'd53479;
   lutrom[1245] = 16'd53508;
   lutrom[1246] = 16'd53537;
   lutrom[1247] = 16'd53566;
   lutrom[1248] = 16'd53595;
   lutrom[1249] = 16'd53624;
   lutrom[1250] = 16'd53653;
   lutrom[1251] = 16'd53682;
   lutrom[1252] = 16'd53710;
   lutrom[1253] = 16'd53739;
   lutrom[1254] = 16'd53768;
   lutrom[1255] = 16'd53797;
   lutrom[1256] = 16'd53825;
   lutrom[1257] = 16'd53854;
   lutrom[1258] = 16'd53883;
   lutrom[1259] = 16'd53911;
   lutrom[1260] = 16'd53940;
   lutrom[1261] = 16'd53968;
   lutrom[1262] = 16'd53997;
   lutrom[1263] = 16'd54025;
   lutrom[1264] = 16'd54054;
   lutrom[1265] = 16'd54082;
   lutrom[1266] = 16'd54110;
   lutrom[1267] = 16'd54139;
   lutrom[1268] = 16'd54167;
   lutrom[1269] = 16'd54195;
   lutrom[1270] = 16'd54224;
   lutrom[1271] = 16'd54252;
   lutrom[1272] = 16'd54280;
   lutrom[1273] = 16'd54308;
   lutrom[1274] = 16'd54336;
   lutrom[1275] = 16'd54364;
   lutrom[1276] = 16'd54392;
   lutrom[1277] = 16'd54420;
   lutrom[1278] = 16'd54448;
   lutrom[1279] = 16'd54476;
   lutrom[1280] = 16'd54504;
   lutrom[1281] = 16'd54532;
   lutrom[1282] = 16'd54560;
   lutrom[1283] = 16'd54588;
   lutrom[1284] = 16'd54616;
   lutrom[1285] = 16'd54643;
   lutrom[1286] = 16'd54671;
   lutrom[1287] = 16'd54699;
   lutrom[1288] = 16'd54727;
   lutrom[1289] = 16'd54754;
   lutrom[1290] = 16'd54782;
   lutrom[1291] = 16'd54809;
   lutrom[1292] = 16'd54837;
   lutrom[1293] = 16'd54864;
   lutrom[1294] = 16'd54892;
   lutrom[1295] = 16'd54919;
   lutrom[1296] = 16'd54947;
   lutrom[1297] = 16'd54974;
   lutrom[1298] = 16'd55001;
   lutrom[1299] = 16'd55029;
   lutrom[1300] = 16'd55056;
   lutrom[1301] = 16'd55083;
   lutrom[1302] = 16'd55111;
   lutrom[1303] = 16'd55138;
   lutrom[1304] = 16'd55165;
   lutrom[1305] = 16'd55192;
   lutrom[1306] = 16'd55219;
   lutrom[1307] = 16'd55246;
   lutrom[1308] = 16'd55273;
   lutrom[1309] = 16'd55300;
   lutrom[1310] = 16'd55327;
   lutrom[1311] = 16'd55354;
   lutrom[1312] = 16'd55381;
   lutrom[1313] = 16'd55408;
   lutrom[1314] = 16'd55435;
   lutrom[1315] = 16'd55461;
   lutrom[1316] = 16'd55488;
   lutrom[1317] = 16'd55515;
   lutrom[1318] = 16'd55542;
   lutrom[1319] = 16'd55568;
   lutrom[1320] = 16'd55595;
   lutrom[1321] = 16'd55621;
   lutrom[1322] = 16'd55648;
   lutrom[1323] = 16'd55675;
   lutrom[1324] = 16'd55701;
   lutrom[1325] = 16'd55728;
   lutrom[1326] = 16'd55754;
   lutrom[1327] = 16'd55780;
   lutrom[1328] = 16'd55807;
   lutrom[1329] = 16'd55833;
   lutrom[1330] = 16'd55859;
   lutrom[1331] = 16'd55886;
   lutrom[1332] = 16'd55912;
   lutrom[1333] = 16'd55938;
   lutrom[1334] = 16'd55964;
   lutrom[1335] = 16'd55990;
   lutrom[1336] = 16'd56017;
   lutrom[1337] = 16'd56043;
   lutrom[1338] = 16'd56069;
   lutrom[1339] = 16'd56095;
   lutrom[1340] = 16'd56121;
   lutrom[1341] = 16'd56147;
   lutrom[1342] = 16'd56172;
   lutrom[1343] = 16'd56198;
   lutrom[1344] = 16'd56224;
   lutrom[1345] = 16'd56250;
   lutrom[1346] = 16'd56276;
   lutrom[1347] = 16'd56301;
   lutrom[1348] = 16'd56327;
   lutrom[1349] = 16'd56353;
   lutrom[1350] = 16'd56379;
   lutrom[1351] = 16'd56404;
   lutrom[1352] = 16'd56430;
   lutrom[1353] = 16'd56455;
   lutrom[1354] = 16'd56481;
   lutrom[1355] = 16'd56506;
   lutrom[1356] = 16'd56532;
   lutrom[1357] = 16'd56557;
   lutrom[1358] = 16'd56582;
   lutrom[1359] = 16'd56608;
   lutrom[1360] = 16'd56633;
   lutrom[1361] = 16'd56658;
   lutrom[1362] = 16'd56684;
   lutrom[1363] = 16'd56709;
   lutrom[1364] = 16'd56734;
   lutrom[1365] = 16'd56759;
   lutrom[1366] = 16'd56784;
   lutrom[1367] = 16'd56809;
   lutrom[1368] = 16'd56834;
   lutrom[1369] = 16'd56859;
   lutrom[1370] = 16'd56884;
   lutrom[1371] = 16'd56909;
   lutrom[1372] = 16'd56934;
   lutrom[1373] = 16'd56959;
   lutrom[1374] = 16'd56984;
   lutrom[1375] = 16'd57009;
   lutrom[1376] = 16'd57034;
   lutrom[1377] = 16'd57058;
   lutrom[1378] = 16'd57083;
   lutrom[1379] = 16'd57108;
   lutrom[1380] = 16'd57132;
   lutrom[1381] = 16'd57157;
   lutrom[1382] = 16'd57181;
   lutrom[1383] = 16'd57206;
   lutrom[1384] = 16'd57231;
   lutrom[1385] = 16'd57255;
   lutrom[1386] = 16'd57279;
   lutrom[1387] = 16'd57304;
   lutrom[1388] = 16'd57328;
   lutrom[1389] = 16'd57353;
   lutrom[1390] = 16'd57377;
   lutrom[1391] = 16'd57401;
   lutrom[1392] = 16'd57425;
   lutrom[1393] = 16'd57450;
   lutrom[1394] = 16'd57474;
   lutrom[1395] = 16'd57498;
   lutrom[1396] = 16'd57522;
   lutrom[1397] = 16'd57546;
   lutrom[1398] = 16'd57570;
   lutrom[1399] = 16'd57594;
   lutrom[1400] = 16'd57618;
   lutrom[1401] = 16'd57642;
   lutrom[1402] = 16'd57666;
   lutrom[1403] = 16'd57690;
   lutrom[1404] = 16'd57714;
   lutrom[1405] = 16'd57737;
   lutrom[1406] = 16'd57761;
   lutrom[1407] = 16'd57785;
   lutrom[1408] = 16'd57809;
   lutrom[1409] = 16'd57832;
   lutrom[1410] = 16'd57856;
   lutrom[1411] = 16'd57879;
   lutrom[1412] = 16'd57903;
   lutrom[1413] = 16'd57927;
   lutrom[1414] = 16'd57950;
   lutrom[1415] = 16'd57973;
   lutrom[1416] = 16'd57997;
   lutrom[1417] = 16'd58020;
   lutrom[1418] = 16'd58044;
   lutrom[1419] = 16'd58067;
   lutrom[1420] = 16'd58090;
   lutrom[1421] = 16'd58113;
   lutrom[1422] = 16'd58137;
   lutrom[1423] = 16'd58160;
   lutrom[1424] = 16'd58183;
   lutrom[1425] = 16'd58206;
   lutrom[1426] = 16'd58229;
   lutrom[1427] = 16'd58252;
   lutrom[1428] = 16'd58275;
   lutrom[1429] = 16'd58298;
   lutrom[1430] = 16'd58321;
   lutrom[1431] = 16'd58344;
   lutrom[1432] = 16'd58367;
   lutrom[1433] = 16'd58390;
   lutrom[1434] = 16'd58413;
   lutrom[1435] = 16'd58435;
   lutrom[1436] = 16'd58458;
   lutrom[1437] = 16'd58481;
   lutrom[1438] = 16'd58504;
   lutrom[1439] = 16'd58526;
   lutrom[1440] = 16'd58549;
   lutrom[1441] = 16'd58571;
   lutrom[1442] = 16'd58594;
   lutrom[1443] = 16'd58616;
   lutrom[1444] = 16'd58639;
   lutrom[1445] = 16'd58661;
   lutrom[1446] = 16'd58684;
   lutrom[1447] = 16'd58706;
   lutrom[1448] = 16'd58728;
   lutrom[1449] = 16'd58751;
   lutrom[1450] = 16'd58773;
   lutrom[1451] = 16'd58795;
   lutrom[1452] = 16'd58817;
   lutrom[1453] = 16'd58839;
   lutrom[1454] = 16'd58862;
   lutrom[1455] = 16'd58884;
   lutrom[1456] = 16'd58906;
   lutrom[1457] = 16'd58928;
   lutrom[1458] = 16'd58950;
   lutrom[1459] = 16'd58972;
   lutrom[1460] = 16'd58993;
   lutrom[1461] = 16'd59015;
   lutrom[1462] = 16'd59037;
   lutrom[1463] = 16'd59059;
   lutrom[1464] = 16'd59081;
   lutrom[1465] = 16'd59103;
   lutrom[1466] = 16'd59124;
   lutrom[1467] = 16'd59146;
   lutrom[1468] = 16'd59168;
   lutrom[1469] = 16'd59189;
   lutrom[1470] = 16'd59211;
   lutrom[1471] = 16'd59232;
   lutrom[1472] = 16'd59254;
   lutrom[1473] = 16'd59275;
   lutrom[1474] = 16'd59297;
   lutrom[1475] = 16'd59318;
   lutrom[1476] = 16'd59339;
   lutrom[1477] = 16'd59361;
   lutrom[1478] = 16'd59382;
   lutrom[1479] = 16'd59403;
   lutrom[1480] = 16'd59424;
   lutrom[1481] = 16'd59446;
   lutrom[1482] = 16'd59467;
   lutrom[1483] = 16'd59488;
   lutrom[1484] = 16'd59509;
   lutrom[1485] = 16'd59530;
   lutrom[1486] = 16'd59551;
   lutrom[1487] = 16'd59572;
   lutrom[1488] = 16'd59593;
   lutrom[1489] = 16'd59614;
   lutrom[1490] = 16'd59635;
   lutrom[1491] = 16'd59655;
   lutrom[1492] = 16'd59676;
   lutrom[1493] = 16'd59697;
   lutrom[1494] = 16'd59718;
   lutrom[1495] = 16'd59738;
   lutrom[1496] = 16'd59759;
   lutrom[1497] = 16'd59780;
   lutrom[1498] = 16'd59800;
   lutrom[1499] = 16'd59821;
   lutrom[1500] = 16'd59841;
   lutrom[1501] = 16'd59862;
   lutrom[1502] = 16'd59882;
   lutrom[1503] = 16'd59903;
   lutrom[1504] = 16'd59923;
   lutrom[1505] = 16'd59943;
   lutrom[1506] = 16'd59964;
   lutrom[1507] = 16'd59984;
   lutrom[1508] = 16'd60004;
   lutrom[1509] = 16'd60024;
   lutrom[1510] = 16'd60044;
   lutrom[1511] = 16'd60065;
   lutrom[1512] = 16'd60085;
   lutrom[1513] = 16'd60105;
   lutrom[1514] = 16'd60125;
   lutrom[1515] = 16'd60145;
   lutrom[1516] = 16'd60165;
   lutrom[1517] = 16'd60185;
   lutrom[1518] = 16'd60204;
   lutrom[1519] = 16'd60224;
   lutrom[1520] = 16'd60244;
   lutrom[1521] = 16'd60264;
   lutrom[1522] = 16'd60284;
   lutrom[1523] = 16'd60303;
   lutrom[1524] = 16'd60323;
   lutrom[1525] = 16'd60343;
   lutrom[1526] = 16'd60362;
   lutrom[1527] = 16'd60382;
   lutrom[1528] = 16'd60401;
   lutrom[1529] = 16'd60421;
   lutrom[1530] = 16'd60440;
   lutrom[1531] = 16'd60460;
   lutrom[1532] = 16'd60479;
   lutrom[1533] = 16'd60498;
   lutrom[1534] = 16'd60518;
   lutrom[1535] = 16'd60537;
   lutrom[1536] = 16'd60556;
   lutrom[1537] = 16'd60575;
   lutrom[1538] = 16'd60594;
   lutrom[1539] = 16'd60614;
   lutrom[1540] = 16'd60633;
   lutrom[1541] = 16'd60652;
   lutrom[1542] = 16'd60671;
   lutrom[1543] = 16'd60690;
   lutrom[1544] = 16'd60709;
   lutrom[1545] = 16'd60728;
   lutrom[1546] = 16'd60746;
   lutrom[1547] = 16'd60765;
   lutrom[1548] = 16'd60784;
   lutrom[1549] = 16'd60803;
   lutrom[1550] = 16'd60822;
   lutrom[1551] = 16'd60840;
   lutrom[1552] = 16'd60859;
   lutrom[1553] = 16'd60878;
   lutrom[1554] = 16'd60896;
   lutrom[1555] = 16'd60915;
   lutrom[1556] = 16'd60933;
   lutrom[1557] = 16'd60952;
   lutrom[1558] = 16'd60970;
   lutrom[1559] = 16'd60989;
   lutrom[1560] = 16'd61007;
   lutrom[1561] = 16'd61025;
   lutrom[1562] = 16'd61044;
   lutrom[1563] = 16'd61062;
   lutrom[1564] = 16'd61080;
   lutrom[1565] = 16'd61098;
   lutrom[1566] = 16'd61117;
   lutrom[1567] = 16'd61135;
   lutrom[1568] = 16'd61153;
   lutrom[1569] = 16'd61171;
   lutrom[1570] = 16'd61189;
   lutrom[1571] = 16'd61207;
   lutrom[1572] = 16'd61225;
   lutrom[1573] = 16'd61243;
   lutrom[1574] = 16'd61261;
   lutrom[1575] = 16'd61278;
   lutrom[1576] = 16'd61296;
   lutrom[1577] = 16'd61314;
   lutrom[1578] = 16'd61332;
   lutrom[1579] = 16'd61349;
   lutrom[1580] = 16'd61367;
   lutrom[1581] = 16'd61385;
   lutrom[1582] = 16'd61402;
   lutrom[1583] = 16'd61420;
   lutrom[1584] = 16'd61437;
   lutrom[1585] = 16'd61455;
   lutrom[1586] = 16'd61472;
   lutrom[1587] = 16'd61490;
   lutrom[1588] = 16'd61507;
   lutrom[1589] = 16'd61524;
   lutrom[1590] = 16'd61542;
   lutrom[1591] = 16'd61559;
   lutrom[1592] = 16'd61576;
   lutrom[1593] = 16'd61593;
   lutrom[1594] = 16'd61610;
   lutrom[1595] = 16'd61628;
   lutrom[1596] = 16'd61645;
   lutrom[1597] = 16'd61662;
   lutrom[1598] = 16'd61679;
   lutrom[1599] = 16'd61696;
   lutrom[1600] = 16'd61713;
   lutrom[1601] = 16'd61729;
   lutrom[1602] = 16'd61746;
   lutrom[1603] = 16'd61763;
   lutrom[1604] = 16'd61780;
   lutrom[1605] = 16'd61797;
   lutrom[1606] = 16'd61813;
   lutrom[1607] = 16'd61830;
   lutrom[1608] = 16'd61847;
   lutrom[1609] = 16'd61863;
   lutrom[1610] = 16'd61880;
   lutrom[1611] = 16'd61896;
   lutrom[1612] = 16'd61913;
   lutrom[1613] = 16'd61929;
   lutrom[1614] = 16'd61946;
   lutrom[1615] = 16'd61962;
   lutrom[1616] = 16'd61979;
   lutrom[1617] = 16'd61995;
   lutrom[1618] = 16'd62011;
   lutrom[1619] = 16'd62027;
   lutrom[1620] = 16'd62044;
   lutrom[1621] = 16'd62060;
   lutrom[1622] = 16'd62076;
   lutrom[1623] = 16'd62092;
   lutrom[1624] = 16'd62108;
   lutrom[1625] = 16'd62124;
   lutrom[1626] = 16'd62140;
   lutrom[1627] = 16'd62156;
   lutrom[1628] = 16'd62172;
   lutrom[1629] = 16'd62188;
   lutrom[1630] = 16'd62204;
   lutrom[1631] = 16'd62219;
   lutrom[1632] = 16'd62235;
   lutrom[1633] = 16'd62251;
   lutrom[1634] = 16'd62267;
   lutrom[1635] = 16'd62282;
   lutrom[1636] = 16'd62298;
   lutrom[1637] = 16'd62313;
   lutrom[1638] = 16'd62329;
   lutrom[1639] = 16'd62345;
   lutrom[1640] = 16'd62360;
   lutrom[1641] = 16'd62375;
   lutrom[1642] = 16'd62391;
   lutrom[1643] = 16'd62406;
   lutrom[1644] = 16'd62422;
   lutrom[1645] = 16'd62437;
   lutrom[1646] = 16'd62452;
   lutrom[1647] = 16'd62467;
   lutrom[1648] = 16'd62482;
   lutrom[1649] = 16'd62498;
   lutrom[1650] = 16'd62513;
   lutrom[1651] = 16'd62528;
   lutrom[1652] = 16'd62543;
   lutrom[1653] = 16'd62558;
   lutrom[1654] = 16'd62573;
   lutrom[1655] = 16'd62588;
   lutrom[1656] = 16'd62603;
   lutrom[1657] = 16'd62617;
   lutrom[1658] = 16'd62632;
   lutrom[1659] = 16'd62647;
   lutrom[1660] = 16'd62662;
   lutrom[1661] = 16'd62676;
   lutrom[1662] = 16'd62691;
   lutrom[1663] = 16'd62706;
   lutrom[1664] = 16'd62720;
   lutrom[1665] = 16'd62735;
   lutrom[1666] = 16'd62749;
   lutrom[1667] = 16'd62764;
   lutrom[1668] = 16'd62778;
   lutrom[1669] = 16'd62793;
   lutrom[1670] = 16'd62807;
   lutrom[1671] = 16'd62821;
   lutrom[1672] = 16'd62836;
   lutrom[1673] = 16'd62850;
   lutrom[1674] = 16'd62864;
   lutrom[1675] = 16'd62878;
   lutrom[1676] = 16'd62893;
   lutrom[1677] = 16'd62907;
   lutrom[1678] = 16'd62921;
   lutrom[1679] = 16'd62935;
   lutrom[1680] = 16'd62949;
   lutrom[1681] = 16'd62963;
   lutrom[1682] = 16'd62977;
   lutrom[1683] = 16'd62991;
   lutrom[1684] = 16'd63004;
   lutrom[1685] = 16'd63018;
   lutrom[1686] = 16'd63032;
   lutrom[1687] = 16'd63046;
   lutrom[1688] = 16'd63059;
   lutrom[1689] = 16'd63073;
   lutrom[1690] = 16'd63087;
   lutrom[1691] = 16'd63100;
   lutrom[1692] = 16'd63114;
   lutrom[1693] = 16'd63127;
   lutrom[1694] = 16'd63141;
   lutrom[1695] = 16'd63154;
   lutrom[1696] = 16'd63168;
   lutrom[1697] = 16'd63181;
   lutrom[1698] = 16'd63194;
   lutrom[1699] = 16'd63208;
   lutrom[1700] = 16'd63221;
   lutrom[1701] = 16'd63234;
   lutrom[1702] = 16'd63247;
   lutrom[1703] = 16'd63261;
   lutrom[1704] = 16'd63274;
   lutrom[1705] = 16'd63287;
   lutrom[1706] = 16'd63300;
   lutrom[1707] = 16'd63313;
   lutrom[1708] = 16'd63326;
   lutrom[1709] = 16'd63339;
   lutrom[1710] = 16'd63352;
   lutrom[1711] = 16'd63364;
   lutrom[1712] = 16'd63377;
   lutrom[1713] = 16'd63390;
   lutrom[1714] = 16'd63403;
   lutrom[1715] = 16'd63415;
   lutrom[1716] = 16'd63428;
   lutrom[1717] = 16'd63441;
   lutrom[1718] = 16'd63453;
   lutrom[1719] = 16'd63466;
   lutrom[1720] = 16'd63478;
   lutrom[1721] = 16'd63491;
   lutrom[1722] = 16'd63503;
   lutrom[1723] = 16'd63516;
   lutrom[1724] = 16'd63528;
   lutrom[1725] = 16'd63540;
   lutrom[1726] = 16'd63553;
   lutrom[1727] = 16'd63565;
   lutrom[1728] = 16'd63577;
   lutrom[1729] = 16'd63589;
   lutrom[1730] = 16'd63601;
   lutrom[1731] = 16'd63614;
   lutrom[1732] = 16'd63626;
   lutrom[1733] = 16'd63638;
   lutrom[1734] = 16'd63650;
   lutrom[1735] = 16'd63662;
   lutrom[1736] = 16'd63673;
   lutrom[1737] = 16'd63685;
   lutrom[1738] = 16'd63697;
   lutrom[1739] = 16'd63709;
   lutrom[1740] = 16'd63721;
   lutrom[1741] = 16'd63732;
   lutrom[1742] = 16'd63744;
   lutrom[1743] = 16'd63756;
   lutrom[1744] = 16'd63767;
   lutrom[1745] = 16'd63779;
   lutrom[1746] = 16'd63791;
   lutrom[1747] = 16'd63802;
   lutrom[1748] = 16'd63814;
   lutrom[1749] = 16'd63825;
   lutrom[1750] = 16'd63836;
   lutrom[1751] = 16'd63848;
   lutrom[1752] = 16'd63859;
   lutrom[1753] = 16'd63870;
   lutrom[1754] = 16'd63881;
   lutrom[1755] = 16'd63893;
   lutrom[1756] = 16'd63904;
   lutrom[1757] = 16'd63915;
   lutrom[1758] = 16'd63926;
   lutrom[1759] = 16'd63937;
   lutrom[1760] = 16'd63948;
   lutrom[1761] = 16'd63959;
   lutrom[1762] = 16'd63970;
   lutrom[1763] = 16'd63981;
   lutrom[1764] = 16'd63992;
   lutrom[1765] = 16'd64003;
   lutrom[1766] = 16'd64013;
   lutrom[1767] = 16'd64024;
   lutrom[1768] = 16'd64035;
   lutrom[1769] = 16'd64046;
   lutrom[1770] = 16'd64056;
   lutrom[1771] = 16'd64067;
   lutrom[1772] = 16'd64077;
   lutrom[1773] = 16'd64088;
   lutrom[1774] = 16'd64098;
   lutrom[1775] = 16'd64109;
   lutrom[1776] = 16'd64119;
   lutrom[1777] = 16'd64130;
   lutrom[1778] = 16'd64140;
   lutrom[1779] = 16'd64150;
   lutrom[1780] = 16'd64160;
   lutrom[1781] = 16'd64171;
   lutrom[1782] = 16'd64181;
   lutrom[1783] = 16'd64191;
   lutrom[1784] = 16'd64201;
   lutrom[1785] = 16'd64211;
   lutrom[1786] = 16'd64221;
   lutrom[1787] = 16'd64231;
   lutrom[1788] = 16'd64241;
   lutrom[1789] = 16'd64251;
   lutrom[1790] = 16'd64261;
   lutrom[1791] = 16'd64271;
   lutrom[1792] = 16'd64281;
   lutrom[1793] = 16'd64290;
   lutrom[1794] = 16'd64300;
   lutrom[1795] = 16'd64310;
   lutrom[1796] = 16'd64320;
   lutrom[1797] = 16'd64329;
   lutrom[1798] = 16'd64339;
   lutrom[1799] = 16'd64348;
   lutrom[1800] = 16'd64358;
   lutrom[1801] = 16'd64367;
   lutrom[1802] = 16'd64377;
   lutrom[1803] = 16'd64386;
   lutrom[1804] = 16'd64395;
   lutrom[1805] = 16'd64405;
   lutrom[1806] = 16'd64414;
   lutrom[1807] = 16'd64423;
   lutrom[1808] = 16'd64432;
   lutrom[1809] = 16'd64442;
   lutrom[1810] = 16'd64451;
   lutrom[1811] = 16'd64460;
   lutrom[1812] = 16'd64469;
   lutrom[1813] = 16'd64478;
   lutrom[1814] = 16'd64487;
   lutrom[1815] = 16'd64496;
   lutrom[1816] = 16'd64505;
   lutrom[1817] = 16'd64514;
   lutrom[1818] = 16'd64522;
   lutrom[1819] = 16'd64531;
   lutrom[1820] = 16'd64540;
   lutrom[1821] = 16'd64549;
   lutrom[1822] = 16'd64557;
   lutrom[1823] = 16'd64566;
   lutrom[1824] = 16'd64574;
   lutrom[1825] = 16'd64583;
   lutrom[1826] = 16'd64592;
   lutrom[1827] = 16'd64600;
   lutrom[1828] = 16'd64608;
   lutrom[1829] = 16'd64617;
   lutrom[1830] = 16'd64625;
   lutrom[1831] = 16'd64634;
   lutrom[1832] = 16'd64642;
   lutrom[1833] = 16'd64650;
   lutrom[1834] = 16'd64658;
   lutrom[1835] = 16'd64666;
   lutrom[1836] = 16'd64675;
   lutrom[1837] = 16'd64683;
   lutrom[1838] = 16'd64691;
   lutrom[1839] = 16'd64699;
   lutrom[1840] = 16'd64707;
   lutrom[1841] = 16'd64715;
   lutrom[1842] = 16'd64723;
   lutrom[1843] = 16'd64731;
   lutrom[1844] = 16'd64738;
   lutrom[1845] = 16'd64746;
   lutrom[1846] = 16'd64754;
   lutrom[1847] = 16'd64762;
   lutrom[1848] = 16'd64769;
   lutrom[1849] = 16'd64777;
   lutrom[1850] = 16'd64785;
   lutrom[1851] = 16'd64792;
   lutrom[1852] = 16'd64800;
   lutrom[1853] = 16'd64807;
   lutrom[1854] = 16'd64815;
   lutrom[1855] = 16'd64822;
   lutrom[1856] = 16'd64829;
   lutrom[1857] = 16'd64837;
   lutrom[1858] = 16'd64844;
   lutrom[1859] = 16'd64851;
   lutrom[1860] = 16'd64858;
   lutrom[1861] = 16'd64866;
   lutrom[1862] = 16'd64873;
   lutrom[1863] = 16'd64880;
   lutrom[1864] = 16'd64887;
   lutrom[1865] = 16'd64894;
   lutrom[1866] = 16'd64901;
   lutrom[1867] = 16'd64908;
   lutrom[1868] = 16'd64915;
   lutrom[1869] = 16'd64922;
   lutrom[1870] = 16'd64929;
   lutrom[1871] = 16'd64935;
   lutrom[1872] = 16'd64942;
   lutrom[1873] = 16'd64949;
   lutrom[1874] = 16'd64956;
   lutrom[1875] = 16'd64962;
   lutrom[1876] = 16'd64969;
   lutrom[1877] = 16'd64975;
   lutrom[1878] = 16'd64982;
   lutrom[1879] = 16'd64988;
   lutrom[1880] = 16'd64995;
   lutrom[1881] = 16'd65001;
   lutrom[1882] = 16'd65008;
   lutrom[1883] = 16'd65014;
   lutrom[1884] = 16'd65020;
   lutrom[1885] = 16'd65027;
   lutrom[1886] = 16'd65033;
   lutrom[1887] = 16'd65039;
   lutrom[1888] = 16'd65045;
   lutrom[1889] = 16'd65051;
   lutrom[1890] = 16'd65057;
   lutrom[1891] = 16'd65063;
   lutrom[1892] = 16'd65069;
   lutrom[1893] = 16'd65075;
   lutrom[1894] = 16'd65081;
   lutrom[1895] = 16'd65087;
   lutrom[1896] = 16'd65093;
   lutrom[1897] = 16'd65099;
   lutrom[1898] = 16'd65105;
   lutrom[1899] = 16'd65110;
   lutrom[1900] = 16'd65116;
   lutrom[1901] = 16'd65122;
   lutrom[1902] = 16'd65127;
   lutrom[1903] = 16'd65133;
   lutrom[1904] = 16'd65138;
   lutrom[1905] = 16'd65144;
   lutrom[1906] = 16'd65149;
   lutrom[1907] = 16'd65155;
   lutrom[1908] = 16'd65160;
   lutrom[1909] = 16'd65166;
   lutrom[1910] = 16'd65171;
   lutrom[1911] = 16'd65176;
   lutrom[1912] = 16'd65181;
   lutrom[1913] = 16'd65187;
   lutrom[1914] = 16'd65192;
   lutrom[1915] = 16'd65197;
   lutrom[1916] = 16'd65202;
   lutrom[1917] = 16'd65207;
   lutrom[1918] = 16'd65212;
   lutrom[1919] = 16'd65217;
   lutrom[1920] = 16'd65222;
   lutrom[1921] = 16'd65227;
   lutrom[1922] = 16'd65232;
   lutrom[1923] = 16'd65236;
   lutrom[1924] = 16'd65241;
   lutrom[1925] = 16'd65246;
   lutrom[1926] = 16'd65251;
   lutrom[1927] = 16'd65255;
   lutrom[1928] = 16'd65260;
   lutrom[1929] = 16'd65265;
   lutrom[1930] = 16'd65269;
   lutrom[1931] = 16'd65274;
   lutrom[1932] = 16'd65278;
   lutrom[1933] = 16'd65282;
   lutrom[1934] = 16'd65287;
   lutrom[1935] = 16'd65291;
   lutrom[1936] = 16'd65295;
   lutrom[1937] = 16'd65300;
   lutrom[1938] = 16'd65304;
   lutrom[1939] = 16'd65308;
   lutrom[1940] = 16'd65312;
   lutrom[1941] = 16'd65316;
   lutrom[1942] = 16'd65321;
   lutrom[1943] = 16'd65325;
   lutrom[1944] = 16'd65329;
   lutrom[1945] = 16'd65333;
   lutrom[1946] = 16'd65337;
   lutrom[1947] = 16'd65340;
   lutrom[1948] = 16'd65344;
   lutrom[1949] = 16'd65348;
   lutrom[1950] = 16'd65352;
   lutrom[1951] = 16'd65356;
   lutrom[1952] = 16'd65359;
   lutrom[1953] = 16'd65363;
   lutrom[1954] = 16'd65367;
   lutrom[1955] = 16'd65370;
   lutrom[1956] = 16'd65374;
   lutrom[1957] = 16'd65377;
   lutrom[1958] = 16'd65381;
   lutrom[1959] = 16'd65384;
   lutrom[1960] = 16'd65387;
   lutrom[1961] = 16'd65391;
   lutrom[1962] = 16'd65394;
   lutrom[1963] = 16'd65397;
   lutrom[1964] = 16'd65401;
   lutrom[1965] = 16'd65404;
   lutrom[1966] = 16'd65407;
   lutrom[1967] = 16'd65410;
   lutrom[1968] = 16'd65413;
   lutrom[1969] = 16'd65416;
   lutrom[1970] = 16'd65419;
   lutrom[1971] = 16'd65422;
   lutrom[1972] = 16'd65425;
   lutrom[1973] = 16'd65428;
   lutrom[1974] = 16'd65431;
   lutrom[1975] = 16'd65434;
   lutrom[1976] = 16'd65436;
   lutrom[1977] = 16'd65439;
   lutrom[1978] = 16'd65442;
   lutrom[1979] = 16'd65445;
   lutrom[1980] = 16'd65447;
   lutrom[1981] = 16'd65450;
   lutrom[1982] = 16'd65452;
   lutrom[1983] = 16'd65455;
   lutrom[1984] = 16'd65457;
   lutrom[1985] = 16'd65460;
   lutrom[1986] = 16'd65462;
   lutrom[1987] = 16'd65464;
   lutrom[1988] = 16'd65467;
   lutrom[1989] = 16'd65469;
   lutrom[1990] = 16'd65471;
   lutrom[1991] = 16'd65473;
   lutrom[1992] = 16'd65476;
   lutrom[1993] = 16'd65478;
   lutrom[1994] = 16'd65480;
   lutrom[1995] = 16'd65482;
   lutrom[1996] = 16'd65484;
   lutrom[1997] = 16'd65486;
   lutrom[1998] = 16'd65488;
   lutrom[1999] = 16'd65490;
   lutrom[2000] = 16'd65492;
   lutrom[2001] = 16'd65493;
   lutrom[2002] = 16'd65495;
   lutrom[2003] = 16'd65497;
   lutrom[2004] = 16'd65499;
   lutrom[2005] = 16'd65500;
   lutrom[2006] = 16'd65502;
   lutrom[2007] = 16'd65503;
   lutrom[2008] = 16'd65505;
   lutrom[2009] = 16'd65506;
   lutrom[2010] = 16'd65508;
   lutrom[2011] = 16'd65509;
   lutrom[2012] = 16'd65511;
   lutrom[2013] = 16'd65512;
   lutrom[2014] = 16'd65513;
   lutrom[2015] = 16'd65515;
   lutrom[2016] = 16'd65516;
   lutrom[2017] = 16'd65517;
   lutrom[2018] = 16'd65518;
   lutrom[2019] = 16'd65519;
   lutrom[2020] = 16'd65520;
   lutrom[2021] = 16'd65521;
   lutrom[2022] = 16'd65522;
   lutrom[2023] = 16'd65523;
   lutrom[2024] = 16'd65524;
   lutrom[2025] = 16'd65525;
   lutrom[2026] = 16'd65526;
   lutrom[2027] = 16'd65527;
   lutrom[2028] = 16'd65528;
   lutrom[2029] = 16'd65528;
   lutrom[2030] = 16'd65529;
   lutrom[2031] = 16'd65530;
   lutrom[2032] = 16'd65530;
   lutrom[2033] = 16'd65531;
   lutrom[2034] = 16'd65531;
   lutrom[2035] = 16'd65532;
   lutrom[2036] = 16'd65532;
   lutrom[2037] = 16'd65533;
   lutrom[2038] = 16'd65533;
   lutrom[2039] = 16'd65534;
   lutrom[2040] = 16'd65534;
   lutrom[2041] = 16'd65534;
   lutrom[2042] = 16'd65534;
   lutrom[2043] = 16'd65535;
   lutrom[2044] = 16'd65535;
   lutrom[2045] = 16'd65535;
   lutrom[2046] = 16'd65535;
   lutrom[2047] = 16'd65535;
end

endmodule
